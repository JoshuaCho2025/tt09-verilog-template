/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_koggestone_adder4 (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

    wire [3:0] a,b;
    wire [3:0] sum;
    wire carry_out;

    assign a = ui_in[3:0];
    assign b = ui_in[7:4];

    wire [3:0] p;
    wire [3:0] q;
    wire [3:0] c;

    assign p = a ^ b;
    assign q = a & b;

    wire g1_1, g1_2, g1_3;
    assign g1_1 = g[1] | (p[1] & g[0]);
    assign g1_2 = g[2] | (p[2] & g[1]);
    assign g1_3 = g[3] | (p[3] & g[2]);

    wire g2_2, g2_3;
    assign g2_2 = g1_2 | (p[2] & g[0]);
    assign g2_3 = g1_3 | (p[3] & g1_1);

    assign c[0] = 0;
    assign c[1] = g[0];
    assign c[2] = g1_1;
    assign c[3] = g2_2;
    assign carry_out = g2_3;

    assign sum = p ^ c;

    assign uo_out[3:0] = sum;
    assign uo_out[4] = carry_out;
    assign uo_out[7:5] = 3'b000;
    assign uio_out = 8'b00000000;
    assign uio_oe = 8'b00000000;
endmodule
  // All output pins must be assigned. If not used, assign to 0.

  // List all unused inputs to prevent warnings
